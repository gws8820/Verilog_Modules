module not_m(A,Y);

input A;
output Y;

nand_m m1(A,A,Y);

endmodule
